









module skid_buffer_tb (
	
);

  // Write your logic here...

endmodule